module XOR2 (y, a, b);
input a, b;
output y;

xor2 x2 (.y(y), .a(a), .b(b));

endmodule

