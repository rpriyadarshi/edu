module AND2 (y, a, b);
input a, b;
output y;

and2 a2 (.y(y), .a(a), .b(b));

endmodule

