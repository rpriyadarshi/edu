module OR2 (y, a, b);
input a, b;
output y;

or o2 (.y(y), .a(a), .b(b));

endmodule

